package baud_rates;

  typedef enum logic [3:0] {
    Br115200,
    Br50,
    Br75,
    Br109_92,
    Br134_51,
    Br150,
    Br300,
    Br600,
    Br1200,
    Br1800,
    Br2400,
    Br3600,
    Br4800,
    Br7200,
    Br9600,
    Br19200
  } baud_rate_t;

endpackage
